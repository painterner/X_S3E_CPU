library verilog;
use verilog.vl_types.all;
entity bus_top is
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        \m0_req_\       : in     vl_logic;
        \m1_req_\       : in     vl_logic;
        \m2_req_\       : in     vl_logic;
        \m3_req_\       : in     vl_logic;
        \m0_grnt_\      : out    vl_logic;
        \m1_grnt_\      : out    vl_logic;
        \m2_grnt_\      : out    vl_logic;
        \m3_grnt_\      : out    vl_logic;
        m0_addr         : in     vl_logic_vector(29 downto 0);
        \m0_as_\        : in     vl_logic;
        m0_rw           : in     vl_logic;
        m0_wr_data      : in     vl_logic_vector(31 downto 0);
        m1_addr         : in     vl_logic_vector(29 downto 0);
        \m1_as_\        : in     vl_logic;
        m1_rw           : in     vl_logic;
        m1_wr_data      : in     vl_logic_vector(31 downto 0);
        m2_addr         : in     vl_logic_vector(29 downto 0);
        \m2_as_\        : in     vl_logic;
        m2_rw           : in     vl_logic;
        m2_wr_data      : in     vl_logic_vector(31 downto 0);
        m3_addr         : in     vl_logic_vector(29 downto 0);
        \m3_as_\        : in     vl_logic;
        m3_rw           : in     vl_logic;
        m3_wr_data      : in     vl_logic_vector(31 downto 0);
        \s0_cs_\        : out    vl_logic;
        \s1_cs_\        : out    vl_logic;
        \s2_cs_\        : out    vl_logic;
        \s3_cs_\        : out    vl_logic;
        \s4_cs_\        : out    vl_logic;
        \s5_cs_\        : out    vl_logic;
        \s6_cs_\        : out    vl_logic;
        \s7_cs_\        : out    vl_logic;
        s_addr          : out    vl_logic_vector(29 downto 0);
        \s_as_\         : out    vl_logic;
        s_rw            : out    vl_logic;
        s_wr_data       : out    vl_logic_vector(31 downto 0);
        s0_rd_data      : in     vl_logic_vector(31 downto 0);
        \s0_rdy_\       : in     vl_logic;
        s1_rd_data      : in     vl_logic_vector(31 downto 0);
        \s1_rdy_\       : in     vl_logic;
        s2_rd_data      : in     vl_logic_vector(31 downto 0);
        \s2_rdy_\       : in     vl_logic;
        s3_rd_data      : in     vl_logic_vector(31 downto 0);
        \s3_rdy_\       : in     vl_logic;
        s4_rd_data      : in     vl_logic_vector(31 downto 0);
        \s4_rdy_\       : in     vl_logic;
        s5_rd_data      : in     vl_logic_vector(31 downto 0);
        \s5_rdy_\       : in     vl_logic;
        s6_rd_data      : in     vl_logic_vector(31 downto 0);
        \s6_rdy_\       : in     vl_logic;
        s7_rd_data      : in     vl_logic_vector(31 downto 0);
        \s7_rdy_\       : in     vl_logic;
        m_rd_data       : out    vl_logic_vector(31 downto 0);
        \m_rdy_\        : out    vl_logic
    );
end bus_top;
