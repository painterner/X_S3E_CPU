
`include "header/firstglobal.h"
`include "header/cpuglobal.h"
`include "header/rom.h"
`include "header/spm.h"
module ctrl(
	input wire							clk,
	input wire							reset,
	
	//***************************************???????
	input wire	[`RegAddrBus]			creg_rd_addr,
	output reg	[`WordDataBus]			creg_rd_data,
	output reg							exe_mode,
	//***************************************??
	input wire	[`CpuIrqBus]			irq,
	output reg							int_detect,
	//***************************************ID/EX??????
	input wire	[`WordAddrBus]			id_pc,
	//***************************************MEM/WB??????
	input wire	[`WordAddrBus]			mem_pc,
	input wire							mem_en,
	input wire							mem_br_flag,
	input wire	[`CtrlOpBus]			mem_ctrl_op,
	input wire	[`RegAddrBus]			mem_dst_addr,
	input wire							mem_gpr_we_,
	input wire	[`IsaExpBus]			mem_exp_code,
	input wire	[`WordDataBus]			mem_out,
	//***************************************??????
	input wire							if_busy,
	input wire							mem_busy,
	input wire							ld_hazard,
	//*************************************** ????
	output wire							if_stall,
	output wire							id_stall,
	output wire							ex_stall,
	output wire							mem_stall,
	//*************************************** ????
	output wire							if_flush,
	output wire							id_flush,
	output wire							ex_flush,
	output wire							mem_flush,
	output reg	[`WordAddrBus]			new_pc

);

	reg									int_en;				//0?????:????
	reg									pre_exe_mode;       //1?????:????
	reg									pre_int_en;         //2?????:????
	reg	[`WordAddrBus]					epc;                //3?????:???????
	reg	[`WordAddrBus]					exp_vector;         //4?????:????
	reg [`IsaExpBus]					exp_code;           //5?????:????
	reg									dly_flag;           //6?????:???????
	reg	[`CpuIrqBus]					mask;               //7?????:????
	reg	[`WordAddrBus]					pre_pc;
	reg									br_flag;
	
	wire	stall				= if_busy|mem_busy;
	assign  if_stall			= stall|ld_hazard;
	assign	id_stall			= stall;
	assign	ex_stall			= stall;
	assign  mem_stall			= stall;
	
	reg		flush;
	assign	if_flush			= flush;
	assign 	id_flush			= flush|ld_hazard;
	assign  ex_flush			= flush;
	assign	mem_flush			= flush;
	
	//******************************************************CPU???????
	always @ *	begin
		new_pc					= `WORD_ADDR_W'H0;
		flush					= `DISABLE;
		if(mem_en == `ENABLE)	
			if(mem_exp_code != `ISA_EXP_NO_EXP)	begin
				new_pc			= exp_vector;
				flush			= `ENABLE;
			end else if(mem_ctrl_op == `CTRL_OP_EXRT)	begin
				new_pc			= epc;
				flush			=`ENABLE;
			end else if(mem_ctrl_op == `CTRL_OP_WRCR)	begin
				new_pc			= mem_pc;
				flush			= `ENABLE;
			end
	end
	
	//******************************************************????
	always @ * 
		if((int_en == `ENABLE) && ((|((~mask) & irq)) == `ENABLE))	
			int_detect			= `ENABLE;
		else
			int_detect			= `DISABLE;
	
	//******************************************************????????
	always @ * 
		case (creg_rd_addr)	
			`CREG_ADDR_STATUS		:																  //   0??????
				creg_rd_data		= {{`WORD_DATA_W-2{1'b0}},int_en,exe_mode};		//??????//  	
			`CREG_ADDR_PRE_STATUS	:                                                                 //   1?????? 
				creg_rd_data		= {{`WORD_DATA_W-2{1'b0}},pre_int_en,pre_exe_mode};                       //   
			`CREG_ADDR_PC			:                                                                 //   2?????? 
				creg_rd_data		= {id_pc,`BYTE_OFFSET_W'H0};                                      //   
			`CREG_ADDR_EPC			:                                                                 //   3?????? 
				creg_rd_data		= {epc,`BYTE_OFFSET_W'H0};                                        //   
			`CREG_ADDR_EXP_VECTOR	:                                                                 //   3?????? 
				creg_rd_data		= {exp_vector,`BYTE_OFFSET_W'H0};                                 //   
			`CREG_ADDR_CAUSE		:                                                                 //   4?????? 
				creg_rd_data		= {{`WORD_DATA_W-1-`ISA_EXP_W{1'H0}},dly_flag,exp_code};          //   
			`CREG_ADDR_INT_MASK		:                                                                 //   5?????? 
				creg_rd_data		= {{`WORD_DATA_W-`CPU_IRQ_CH{1'B0}},mask};                        //   
			`CREG_ADDR_IRQ			:                                                                 //   6?????? 
				creg_rd_data		= {{`WORD_DATA_W-`CPU_IRQ_CH{1'B0}},irq};                         //   
			`CREG_ADDR_ROM_SIZE		:                                                                 //   7?????? 
				creg_rd_data		= $unsigned(`ROM_SIZE);                                           //
			`CREG_ADDR_SPM_SIZE		:                                                                 //  29?????? 
				creg_rd_data		= $unsigned(`SPM_SIZE);                                           //
			`CREG_ADDR_CPU_INFO		:                                                                    //  30? register
				creg_rd_data		= {`RELEASE_YEAR,`RELEASE_MONTH,`RELEASE_VERSION,`RELEASE_REVISION}; //
			default					:                                                                    //  31? register
				creg_rd_data		= `WORD_DATA_W'H0;                                                   //
		endcase

	//******************************************************CPU???
	always @(posedge clk or `RESET_EDGE reset)	
		if(reset == `RESET_ENABLE)	begin
			exe_mode				<= #1 `CPU_KERNEL_MODE;
			int_en					<= #1 `DISABLE;
			pre_exe_mode			<= #1 `CPU_KERNEL_MODE;
			pre_int_en				<= #1 `DISABLE;
			exp_code				<= #1 `ISA_EXP_NO_EXP;
			mask					<= #1 {`CPU_IRQ_CH{`ENABLE}};
			dly_flag				<= #1 `DISABLE;
			epc						<= #1 `WORD_ADDR_W'H0;
			exp_vector				<= #1 `WORD_ADDR_W'H0;
			pre_pc					<= #1 `WORD_ADDR_W'H0;
			br_flag					<= #1 `DISABLE;
		end else
			if((mem_en == `ENABLE) && (stall == `DISABLE))	begin				//pc?????????
				pre_pc				<= #1 mem_pc;
				br_flag				<= #1 mem_br_flag;
				if(mem_exp_code != `ISA_EXP_NO_EXP)	begin					//????
					exe_mode				<= #1 `CPU_KERNEL_MODE;
			        int_en					<= #1 `DISABLE;
			        pre_exe_mode			<= #1 exe_mode;
			        pre_int_en				<= #1 int_en;
			        exp_code				<= #1 mem_exp_code;
			        dly_flag				<= #1 br_flag;
			        epc						<= #1 pre_pc;
			    end else if(mem_ctrl_op == `CTRL_OP_EXRT)	begin			//exrt??
			    	exe_mode				<= #1 pre_exe_mode;
			    	int_en					<= #1 pre_int_en;
			    end else if(mem_ctrl_op == `CTRL_OP_WRCR)				//wrcr??
			    	case(mem_dst_addr)
			    		`CREG_ADDR_STATUS		:	begin								//0??????
			    			exe_mode		<= #1 mem_out[`CregExeModeLoc];
			    			int_en			<= #1 mem_out[`CregIntEnableLoc];
			    		end
			    		`CREG_ADDR_PRE_STATUS		:	begin								//1??????
			    			pre_exe_mode	<= #1 mem_out[`CregExeModeLoc];    
			    			pre_int_en		<= #1 mem_out[`CregIntEnableLoc]; 
			    		end
			    		`CREG_ADDR_EPC			:										//3??????
			    			epc				<= #1 mem_out[`WordAddrLoc];
			    		`CREG_ADDR_EXP_VECTOR	:										//4??????
			    			exp_vector		<= #1 mem_out[`WordAddrLoc]; 
			    		`CREG_ADDR_CAUSE		: begin										//5??????
			    			dly_flag		<= #1 mem_out[`CregDlyFlagLoc];
			    			exp_code		<= #1 mem_out[`CregExpCodeLoc];
			    			end
			    		`CREG_ADDR_INT_MASK	 	:										//6??????
			    			mask			<= #1 mem_out[`CPU_IRQ_CH-1:0];
			    	endcase
			end
					
endmodule		
			    	 
			    			
			   
			    	
					
			
				
				
			
		
		
			
			
	
	
	
