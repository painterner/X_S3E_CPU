`include "header/firstglobal.h"              
`include "header/cpuglobal.h" 

`include "CPU/EX/alu.v"
`include "CPU/EX/ex_reg.v"               
module ex_top(
	input wire							clk   		   ,
    input wire							reset          ,
                                                       
	input wire	[`WordDataBus]				in_0       ,
  	input wire	[`WordDataBus]				in_1       ,
    input wire	[`AluOpBus]					op         ,
                                                       
    //*****************************????            
    input wire							stall          ,
    input wire							flush          ,
    input wire							int_detect	   , 			//????
    //*****************************ID/EX??????   
    input wire	[`WordAddrBus]			id_pc          ,
    input wire							id_en          ,
    input wire							id_br_flag     ,
    input wire	[`MemOpBus]				id_mem_op      ,
    input wire	[`WordDataBus]			id_mem_wr_data ,
    input wire	[`CtrlOpBus ]			id_ctrl_op     ,
    input wire	[`RegAddrBus]			id_dst_addr    ,
    input wire							id_gpr_we_     ,
    input wire	[`IsaExpBus]			id_exp_code    ,
    //*****************************EX/MEM??????  
    output wire	[`WordAddrBus]			ex_pc          ,
    output wire							ex_en          ,
    output wire							ex_br_flag     ,
    output wire	[`MemOpBus]				ex_mem_op      ,
    output wire	[`WordDataBus]			ex_mem_wr_data ,
    output wire	[`CtrlOpBus]			ex_ctrl_op     ,
    output wire	[`RegAddrBus]			ex_dst_addr    ,
    output wire							ex_gpr_we_     ,
    output wire	[`IsaExpBus]			ex_exp_code    ,
    output wire	[`WordDataBus]			ex_out     	   ,
    
    //*****************************************************???**********************//
    output wire	[`WordDataBus]			fwd_data		    			//????
 
 );
 
 	   wire	[`WordDataBus]				out ; 
	   wire								of  ; 
	   assign fwd_data			= out;

 	alu alu(
 	   		.in_0   				(in_0)			,
 	   		.in_1                   (in_1)          ,
 	   		.op                     (op  )          ,
			.out  					(out)           ,
 			.of   					(of)            


 	); 
 	
 	ex_reg ex_reg(
 			.clk					   (clk				  )				,
 			.reset					   (reset			  )				,
 			.stall                     (  stall           ) 			,
 	        .flush                     (  flush           )             ,
 	        .int_detect			       (  int_detect	  )              ,
 	        .id_pc                     (  id_pc           )             ,
 	        .id_en                     (  id_en           )             ,
 	        .id_br_flag                (  id_br_flag      )             ,
 	        .id_mem_op                 (  id_mem_op       )             ,
 	        .id_mem_wr_data            (  id_mem_wr_data  )             ,
 	        .id_ctrl_op                (  id_ctrl_op      )             ,
 	        .id_dst_addr               (  id_dst_addr     )             ,
 	        .id_gpr_we_                (  id_gpr_we_      )             ,
 	        .id_exp_code               (  id_exp_code     )             ,   
 	        .ex_pc                     (  ex_pc           )             ,
 	        .ex_en                     (  ex_en           )             ,
 	        .ex_br_flag                (  ex_br_flag      )             ,
 	        .ex_mem_op                 (  ex_mem_op       )             ,
 	        .ex_mem_wr_data            (  ex_mem_wr_data  )             ,
 	        .ex_ctrl_op                (  ex_ctrl_op      )             ,
 	        .ex_dst_addr               (  ex_dst_addr     )             ,
 	        .ex_gpr_we_                (  ex_gpr_we_      )             ,
 	        .ex_exp_code               (  ex_exp_code     )             ,
 	        .ex_out                    (  ex_out          )             ,
 	        .alu_out				   (	 out		  )             ,
 	        .alu_of      			   (	 of		   	  )              
 	 	
 	) ;

endmodule                                                 
   
   